library verilog;
use verilog.vl_types.all;
entity Top_sv_unit is
end Top_sv_unit;
