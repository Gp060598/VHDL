library verilog;
use verilog.vl_types.all;
entity test_config_reg is
end test_config_reg;
